library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity rom_c64_kernal is
	port (
		clk: in std_logic;
		addr: in unsigned(12 downto 0);
		do: out unsigned(7 downto 0)
	);
end entity;

architecture Behavioral of rom_c64_kernal is
	type romDef is array(0 to  8191) of unsigned(7 downto 0);
	constant romData: romDef := (
		X"85", X"56", X"20", X"0F", X"BC", X"A5", X"61", X"C9", X"88", X"90", X"03", X"20", X"D4", X"BA", X"20", X"CC", 
		X"BC", X"A5", X"07", X"18", X"69", X"81", X"F0", X"F3", X"38", X"E9", X"01", X"48", X"A2", X"05", X"B5", X"69", 
		X"B4", X"61", X"95", X"61", X"94", X"69", X"CA", X"10", X"F5", X"A5", X"56", X"85", X"70", X"20", X"53", X"B8", 
		X"20", X"B4", X"BF", X"A9", X"C4", X"A0", X"BF", X"20", X"59", X"E0", X"A9", X"00", X"85", X"6F", X"68", X"20", 
		X"B9", X"BA", X"60", X"85", X"71", X"84", X"72", X"20", X"CA", X"BB", X"A9", X"57", X"20", X"28", X"BA", X"20", 
		X"5D", X"E0", X"A9", X"57", X"A0", X"00", X"4C", X"28", X"BA", X"85", X"71", X"84", X"72", X"20", X"C7", X"BB", 
		X"B1", X"71", X"85", X"67", X"A4", X"71", X"C8", X"98", X"D0", X"02", X"E6", X"72", X"85", X"71", X"A4", X"72", 
		X"20", X"28", X"BA", X"A5", X"71", X"A4", X"72", X"18", X"69", X"05", X"90", X"01", X"C8", X"85", X"71", X"84", 
		X"72", X"20", X"67", X"B8", X"A9", X"5C", X"A0", X"00", X"C6", X"67", X"D0", X"E4", X"60", X"98", X"35", X"44", 
		X"7A", X"00", X"68", X"28", X"B1", X"46", X"00", X"20", X"2B", X"BC", X"30", X"37", X"D0", X"20", X"20", X"F3", 
		X"FF", X"86", X"22", X"84", X"23", X"A0", X"04", X"B1", X"22", X"85", X"62", X"C8", X"B1", X"22", X"85", X"64", 
		X"A0", X"08", X"B1", X"22", X"85", X"63", X"C8", X"B1", X"22", X"85", X"65", X"4C", X"E3", X"E0", X"A9", X"8B", 
		X"A0", X"00", X"20", X"A2", X"BB", X"A9", X"8D", X"A0", X"E0", X"20", X"28", X"BA", X"A9", X"92", X"A0", X"E0", 
		X"20", X"67", X"B8", X"A6", X"65", X"A5", X"62", X"85", X"65", X"86", X"62", X"A6", X"63", X"A5", X"64", X"85", 
		X"63", X"86", X"64", X"A9", X"00", X"85", X"66", X"A5", X"61", X"85", X"70", X"A9", X"80", X"85", X"61", X"20", 
		X"D7", X"B8", X"A2", X"8B", X"A0", X"00", X"4C", X"D4", X"BB", X"C9", X"F0", X"D0", X"07", X"84", X"38", X"86", 
		X"37", X"4C", X"63", X"A6", X"AA", X"D0", X"02", X"A2", X"1E", X"4C", X"37", X"A4", X"20", X"D2", X"FF", X"B0", 
		X"E8", X"60", X"20", X"CF", X"FF", X"B0", X"E2", X"60", X"20", X"AD", X"E4", X"B0", X"DC", X"60", X"20", X"C6", 
		X"FF", X"B0", X"D6", X"60", X"20", X"E4", X"FF", X"B0", X"D0", X"60", X"20", X"8A", X"AD", X"20", X"F7", X"B7", 
		X"A9", X"E1", X"48", X"A9", X"46", X"48", X"AD", X"0F", X"03", X"48", X"AD", X"0C", X"03", X"AE", X"0D", X"03", 
		X"AC", X"0E", X"03", X"28", X"6C", X"14", X"00", X"08", X"8D", X"0C", X"03", X"8E", X"0D", X"03", X"8C", X"0E", 
		X"03", X"68", X"8D", X"0F", X"03", X"60", X"20", X"D4", X"E1", X"A6", X"2D", X"A4", X"2E", X"A9", X"2B", X"20", 
		X"D8", X"FF", X"B0", X"95", X"60", X"A9", X"01", X"2C", X"A9", X"00", X"85", X"0A", X"20", X"D4", X"E1", X"A5", 
		X"0A", X"A6", X"2B", X"A4", X"2C", X"20", X"D5", X"FF", X"B0", X"57", X"A5", X"0A", X"F0", X"17", X"A2", X"1C", 
		X"20", X"B7", X"FF", X"29", X"10", X"D0", X"17", X"A5", X"7A", X"C9", X"02", X"F0", X"07", X"A9", X"64", X"A0", 
		X"A3", X"4C", X"1E", X"AB", X"60", X"20", X"B7", X"FF", X"29", X"BF", X"F0", X"05", X"A2", X"1D", X"4C", X"37", 
		X"A4", X"A5", X"7B", X"C9", X"02", X"D0", X"0E", X"86", X"2D", X"84", X"2E", X"A9", X"76", X"A0", X"A3", X"20", 
		X"1E", X"AB", X"4C", X"2A", X"A5", X"20", X"8E", X"A6", X"20", X"33", X"A5", X"4C", X"77", X"A6", X"20", X"19", 
		X"E2", X"20", X"C0", X"FF", X"B0", X"0B", X"60", X"20", X"19", X"E2", X"A5", X"49", X"20", X"C3", X"FF", X"90", 
		X"C3", X"4C", X"F9", X"E0", X"A9", X"00", X"20", X"BD", X"FF", X"A2", X"01", X"A0", X"00", X"20", X"BA", X"FF", 
		X"20", X"06", X"E2", X"20", X"57", X"E2", X"20", X"06", X"E2", X"20", X"00", X"E2", X"A0", X"00", X"86", X"49", 
		X"20", X"BA", X"FF", X"20", X"06", X"E2", X"20", X"00", X"E2", X"8A", X"A8", X"A6", X"49", X"4C", X"BA", X"FF", 
		X"20", X"0E", X"E2", X"4C", X"9E", X"B7", X"20", X"79", X"00", X"D0", X"02", X"68", X"68", X"60", X"20", X"FD", 
		X"AE", X"20", X"79", X"00", X"D0", X"F7", X"4C", X"08", X"AF", X"A9", X"00", X"20", X"BD", X"FF", X"20", X"11", 
		X"E2", X"20", X"9E", X"B7", X"86", X"49", X"8A", X"A2", X"01", X"A0", X"00", X"20", X"BA", X"FF", X"20", X"06", 
		X"E2", X"20", X"00", X"E2", X"86", X"4A", X"A0", X"00", X"A5", X"49", X"E0", X"03", X"90", X"01", X"88", X"20", 
		X"BA", X"FF", X"20", X"06", X"E2", X"20", X"00", X"E2", X"8A", X"A8", X"A6", X"4A", X"A5", X"49", X"20", X"BA", 
		X"FF", X"20", X"06", X"E2", X"20", X"0E", X"E2", X"20", X"9E", X"AD", X"20", X"A3", X"B6", X"A6", X"22", X"A4", 
		X"23", X"4C", X"BD", X"FF", X"A9", X"E0", X"A0", X"E2", X"20", X"67", X"B8", X"20", X"0C", X"BC", X"A9", X"E5", 
		X"A0", X"E2", X"A6", X"6E", X"20", X"07", X"BB", X"20", X"0C", X"BC", X"20", X"CC", X"BC", X"A9", X"00", X"85", 
		X"6F", X"20", X"53", X"B8", X"A9", X"EA", X"A0", X"E2", X"20", X"50", X"B8", X"A5", X"66", X"48", X"10", X"0D", 
		X"20", X"49", X"B8", X"A5", X"66", X"30", X"09", X"A5", X"12", X"49", X"FF", X"85", X"12", X"20", X"B4", X"BF", 
		X"A9", X"EA", X"A0", X"E2", X"20", X"67", X"B8", X"68", X"10", X"03", X"20", X"B4", X"BF", X"A9", X"EF", X"A0", 
		X"E2", X"4C", X"43", X"E0", X"20", X"CA", X"BB", X"A9", X"00", X"85", X"12", X"20", X"6B", X"E2", X"A2", X"4E", 
		X"A0", X"00", X"20", X"F6", X"E0", X"A9", X"57", X"A0", X"00", X"20", X"A2", X"BB", X"A9", X"00", X"85", X"66", 
		X"A5", X"12", X"20", X"DC", X"E2", X"A9", X"4E", X"A0", X"00", X"4C", X"0F", X"BB", X"48", X"4C", X"9D", X"E2", 
		X"81", X"49", X"0F", X"DA", X"A2", X"83", X"49", X"0F", X"DA", X"A2", X"7F", X"00", X"00", X"00", X"00", X"05", 
		X"84", X"E6", X"1A", X"2D", X"1B", X"86", X"28", X"07", X"FB", X"F8", X"87", X"99", X"68", X"89", X"01", X"87", 
		X"23", X"35", X"DF", X"E1", X"86", X"A5", X"5D", X"E7", X"28", X"83", X"49", X"0F", X"DA", X"A2", X"A5", X"66", 
		X"48", X"10", X"03", X"20", X"B4", X"BF", X"A5", X"61", X"48", X"C9", X"81", X"90", X"07", X"A9", X"BC", X"A0", 
		X"B9", X"20", X"0F", X"BB", X"A9", X"3E", X"A0", X"E3", X"20", X"43", X"E0", X"68", X"C9", X"81", X"90", X"07", 
		X"A9", X"E0", X"A0", X"E2", X"20", X"50", X"B8", X"68", X"10", X"03", X"4C", X"B4", X"BF", X"60", X"0B", X"76", 
		X"B3", X"83", X"BD", X"D3", X"79", X"1E", X"F4", X"A6", X"F5", X"7B", X"83", X"FC", X"B0", X"10", X"7C", X"0C", 
		X"1F", X"67", X"CA", X"7C", X"DE", X"53", X"CB", X"C1", X"7D", X"14", X"64", X"70", X"4C", X"7D", X"B7", X"EA", 
		X"51", X"7A", X"7D", X"63", X"30", X"88", X"7E", X"7E", X"92", X"44", X"99", X"3A", X"7E", X"4C", X"CC", X"91", 
		X"C7", X"7F", X"AA", X"AA", X"AA", X"13", X"81", X"00", X"00", X"00", X"00", X"20", X"CC", X"FF", X"A9", X"00", 
		X"85", X"13", X"20", X"7A", X"A6", X"58", X"A2", X"80", X"6C", X"00", X"03", X"8A", X"30", X"03", X"4C", X"3A", 
		X"A4", X"4C", X"74", X"A4", X"20", X"53", X"E4", X"20", X"BF", X"E3", X"20", X"22", X"E4", X"A2", X"FB", X"9A", 
		X"D0", X"E4", X"E6", X"7A", X"D0", X"02", X"E6", X"7B", X"AD", X"60", X"EA", X"C9", X"3A", X"B0", X"0A", X"C9", 
		X"20", X"F0", X"EF", X"38", X"E9", X"30", X"38", X"E9", X"D0", X"60", X"80", X"4F", X"C7", X"52", X"58", X"A9", 
		X"4C", X"85", X"54", X"8D", X"10", X"03", X"A9", X"48", X"A0", X"B2", X"8D", X"11", X"03", X"8C", X"12", X"03", 
		X"A9", X"91", X"A0", X"B3", X"85", X"05", X"84", X"06", X"A9", X"AA", X"A0", X"B1", X"85", X"03", X"84", X"04", 
		X"A2", X"1C", X"BD", X"A2", X"E3", X"95", X"73", X"CA", X"10", X"F8", X"A9", X"03", X"85", X"53", X"A9", X"00", 
		X"85", X"68", X"85", X"13", X"85", X"18", X"A2", X"01", X"8E", X"FD", X"01", X"8E", X"FC", X"01", X"A2", X"19", 
		X"86", X"16", X"38", X"20", X"9C", X"FF", X"86", X"2B", X"84", X"2C", X"38", X"20", X"99", X"FF", X"86", X"37", 
		X"84", X"38", X"86", X"33", X"84", X"34", X"A0", X"00", X"98", X"91", X"2B", X"E6", X"2B", X"D0", X"02", X"E6", 
		X"2C", X"60", X"A5", X"2B", X"A4", X"2C", X"20", X"08", X"A4", X"A9", X"73", X"A0", X"E4", X"20", X"1E", X"AB", 
		X"A5", X"37", X"38", X"E5", X"2B", X"AA", X"A5", X"38", X"E5", X"2C", X"20", X"CD", X"BD", X"A9", X"60", X"A0", 
		X"E4", X"20", X"1E", X"AB", X"4C", X"44", X"A6", X"8B", X"E3", X"83", X"A4", X"7C", X"A5", X"1A", X"A7", X"E4", 
		X"A7", X"86", X"AE", X"A2", X"0B", X"BD", X"47", X"E4", X"9D", X"00", X"03", X"CA", X"10", X"F7", X"60", X"00", 
		X"20", X"42", X"41", X"53", X"49", X"43", X"20", X"42", X"59", X"54", X"45", X"53", X"20", X"46", X"52", X"45", 
		X"45", X"0D", X"00", X"93", X"0D", X"20", X"20", X"20", X"20", X"2A", X"2A", X"2A", X"2A", X"20", X"43", X"4F", 
		X"4D", X"4D", X"4F", X"44", X"4F", X"52", X"45", X"20", X"36", X"34", X"20", X"42", X"41", X"53", X"49", X"43", 
		X"20", X"56", X"32", X"20", X"2A", X"2A", X"2A", X"2A", X"0D", X"0D", X"20", X"36", X"34", X"4B", X"20", X"52", 
		X"41", X"4D", X"20", X"53", X"59", X"53", X"54", X"45", X"4D", X"20", X"20", X"00", X"81", X"48", X"20", X"C9", 
		X"FF", X"AA", X"68", X"90", X"01", X"8A", X"60", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", 
		X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", X"AA", 
		X"AA", X"AA", X"AA", X"85", X"A9", X"A9", X"01", X"85", X"AB", X"60", X"AD", X"86", X"02", X"91", X"F3", X"60", 
		X"69", X"02", X"A4", X"91", X"C8", X"D0", X"04", X"C5", X"A1", X"D0", X"F7", X"60", X"19", X"26", X"44", X"19", 
		X"1A", X"11", X"E8", X"0D", X"70", X"0C", X"06", X"06", X"D1", X"02", X"37", X"01", X"AE", X"00", X"69", X"00", 
		X"A2", X"00", X"A0", X"DC", X"60", X"A2", X"28", X"A0", X"19", X"60", X"B0", X"07", X"86", X"D6", X"84", X"D3", 
		X"20", X"6C", X"E5", X"A6", X"D6", X"A4", X"D3", X"60", X"20", X"A0", X"E5", X"A9", X"00", X"8D", X"91", X"02", 
		X"85", X"CF", X"A9", X"48", X"8D", X"8F", X"02", X"A9", X"EB", X"8D", X"90", X"02", X"A9", X"0A", X"8D", X"89", 
		X"02", X"8D", X"8C", X"02", X"A9", X"0E", X"8D", X"86", X"02", X"A9", X"04", X"8D", X"8B", X"02", X"A9", X"0C", 
		X"85", X"CD", X"85", X"CC", X"AD", X"88", X"02", X"09", X"80", X"A8", X"A9", X"00", X"AA", X"94", X"D9", X"18", 
		X"69", X"28", X"90", X"01", X"C8", X"E8", X"E0", X"1A", X"D0", X"F3", X"A9", X"FF", X"95", X"D9", X"A2", X"18", 
		X"20", X"FF", X"E9", X"CA", X"10", X"FA", X"A0", X"00", X"84", X"D3", X"84", X"D6", X"A6", X"D6", X"A5", X"D3", 
		X"B4", X"D9", X"30", X"08", X"18", X"69", X"28", X"85", X"D3", X"CA", X"10", X"F4", X"20", X"F0", X"E9", X"A9", 
		X"27", X"E8", X"B4", X"D9", X"30", X"06", X"18", X"69", X"28", X"E8", X"10", X"F6", X"85", X"D5", X"4C", X"24", 
		X"EA", X"E4", X"C9", X"F0", X"03", X"4C", X"ED", X"E6", X"60", X"EA", X"20", X"A0", X"E5", X"4C", X"66", X"E5", 
		X"A9", X"03", X"85", X"9A", X"A9", X"00", X"85", X"99", X"A2", X"2F", X"BD", X"B8", X"EC", X"9D", X"FF", X"CF", 
		X"CA", X"D0", X"F7", X"60", X"AC", X"77", X"02", X"A2", X"00", X"BD", X"78", X"02", X"9D", X"77", X"02", X"E8", 
		X"E4", X"C6", X"D0", X"F5", X"C6", X"C6", X"98", X"58", X"18", X"60", X"20", X"16", X"E7", X"A5", X"C6", X"85", 
		X"CC", X"8D", X"92", X"02", X"F0", X"F7", X"78", X"A5", X"CF", X"F0", X"0C", X"A5", X"CE", X"AE", X"87", X"02", 
		X"A0", X"00", X"84", X"CF", X"20", X"13", X"EA", X"20", X"B4", X"E5", X"C9", X"83", X"D0", X"10", X"A2", X"09", 
		X"78", X"86", X"C6", X"BD", X"E6", X"EC", X"9D", X"76", X"02", X"CA", X"D0", X"F7", X"F0", X"CF", X"C9", X"0D", 
		X"D0", X"C8", X"A4", X"D5", X"84", X"D0", X"B1", X"D1", X"C9", X"20", X"D0", X"03", X"88", X"D0", X"F7", X"C8", 
		X"84", X"C8", X"A0", X"00", X"8C", X"92", X"02", X"84", X"D3", X"84", X"D4", X"A5", X"C9", X"30", X"1B", X"A6", 
		X"D6", X"20", X"91", X"E5", X"E4", X"C9", X"D0", X"12", X"A5", X"CA", X"85", X"D3", X"C5", X"C8", X"90", X"0A", 
		X"B0", X"2B", X"98", X"48", X"8A", X"48", X"A5", X"D0", X"F0", X"93", X"A4", X"D3", X"B1", X"D1", X"85", X"D7", 
		X"29", X"3F", X"06", X"D7", X"24", X"D7", X"10", X"02", X"09", X"80", X"90", X"04", X"A6", X"D4", X"D0", X"04", 
		X"70", X"02", X"09", X"40", X"E6", X"D3", X"20", X"84", X"E6", X"C4", X"C8", X"D0", X"17", X"A9", X"00", X"85", 
		X"D0", X"A9", X"0D", X"A6", X"99", X"E0", X"03", X"F0", X"06", X"A6", X"9A", X"E0", X"03", X"F0", X"03", X"20", 
		X"16", X"E7", X"A9", X"0D", X"85", X"D7", X"68", X"AA", X"68", X"A8", X"A5", X"D7", X"C9", X"DE", X"D0", X"02", 
		X"A9", X"FF", X"18", X"60", X"C9", X"22", X"D0", X"08", X"A5", X"D4", X"49", X"01", X"85", X"D4", X"A9", X"22", 
		X"60", X"09", X"40", X"A6", X"C7", X"F0", X"02", X"09", X"80", X"A6", X"D8", X"F0", X"02", X"C6", X"D8", X"AE", 
		X"86", X"02", X"20", X"13", X"EA", X"20", X"B6", X"E6", X"68", X"A8", X"A5", X"D8", X"F0", X"02", X"46", X"D4", 
		X"68", X"AA", X"68", X"18", X"58", X"60", X"20", X"B3", X"E8", X"E6", X"D3", X"A5", X"D5", X"C5", X"D3", X"B0", 
		X"3F", X"C9", X"4F", X"F0", X"32", X"AD", X"92", X"02", X"F0", X"03", X"4C", X"67", X"E9", X"A6", X"D6", X"E0", 
		X"19", X"90", X"07", X"20", X"EA", X"E8", X"C6", X"D6", X"A6", X"D6", X"16", X"D9", X"56", X"D9", X"E8", X"B5", 
		X"D9", X"09", X"80", X"95", X"D9", X"CA", X"A5", X"D5", X"18", X"69", X"28", X"85", X"D5", X"B5", X"D9", X"30", 
		X"03", X"CA", X"D0", X"F9", X"4C", X"F0", X"E9", X"C6", X"D6", X"20", X"7C", X"E8", X"A9", X"00", X"85", X"D3", 
		X"60", X"A6", X"D6", X"D0", X"06", X"86", X"D3", X"68", X"68", X"D0", X"9D", X"CA", X"86", X"D6", X"20", X"6C", 
		X"E5", X"A4", X"D5", X"84", X"D3", X"60", X"48", X"85", X"D7", X"8A", X"48", X"98", X"48", X"A9", X"00", X"85", 
		X"D0", X"A4", X"D3", X"A5", X"D7", X"10", X"03", X"4C", X"D4", X"E7", X"C9", X"0D", X"D0", X"03", X"4C", X"91", 
		X"E8", X"C9", X"20", X"90", X"10", X"C9", X"60", X"90", X"04", X"29", X"DF", X"D0", X"02", X"29", X"3F", X"20", 
		X"84", X"E6", X"4C", X"93", X"E6", X"A6", X"D8", X"F0", X"03", X"4C", X"97", X"E6", X"C9", X"14", X"D0", X"2E", 
		X"98", X"D0", X"06", X"20", X"01", X"E7", X"4C", X"73", X"E7", X"20", X"A1", X"E8", X"88", X"84", X"D3", X"20", 
		X"24", X"EA", X"C8", X"B1", X"D1", X"88", X"91", X"D1", X"C8", X"B1", X"F3", X"88", X"91", X"F3", X"C8", X"C4", 
		X"D5", X"D0", X"EF", X"A9", X"20", X"91", X"D1", X"AD", X"86", X"02", X"91", X"F3", X"10", X"4D", X"A6", X"D4", 
		X"F0", X"03", X"4C", X"97", X"E6", X"C9", X"12", X"D0", X"02", X"85", X"C7", X"C9", X"13", X"D0", X"03", X"20", 
		X"66", X"E5", X"C9", X"1D", X"D0", X"17", X"C8", X"20", X"B3", X"E8", X"84", X"D3", X"88", X"C4", X"D5", X"90", 
		X"09", X"C6", X"D6", X"20", X"7C", X"E8", X"A0", X"00", X"84", X"D3", X"4C", X"A8", X"E6", X"C9", X"11", X"D0", 
		X"1D", X"18", X"98", X"69", X"28", X"A8", X"E6", X"D6", X"C5", X"D5", X"90", X"EC", X"F0", X"EA", X"C6", X"D6", 
		X"E9", X"28", X"90", X"04", X"85", X"D3", X"D0", X"F8", X"20", X"7C", X"E8", X"4C", X"A8", X"E6", X"20", X"CB", 
		X"E8", X"4C", X"44", X"EC", X"29", X"7F", X"C9", X"7F", X"D0", X"02", X"A9", X"5E", X"C9", X"20", X"90", X"03", 
		X"4C", X"91", X"E6", X"C9", X"0D", X"D0", X"03", X"4C", X"91", X"E8", X"A6", X"D4", X"D0", X"3F", X"C9", X"14", 
		X"D0", X"37", X"A4", X"D5", X"B1", X"D1", X"C9", X"20", X"D0", X"04", X"C4", X"D3", X"D0", X"07", X"C0", X"4F", 
		X"F0", X"24", X"20", X"65", X"E9", X"A4", X"D5", X"20", X"24", X"EA", X"88", X"B1", X"D1", X"C8", X"91", X"D1", 
		X"88", X"B1", X"F3", X"C8", X"91", X"F3", X"88", X"C4", X"D3", X"D0", X"EF", X"A9", X"20", X"91", X"D1", X"AD", 
		X"86", X"02", X"91", X"F3", X"E6", X"D8", X"4C", X"A8", X"E6", X"A6", X"D8", X"F0", X"05", X"09", X"40", X"4C", 
		X"97", X"E6", X"C9", X"11", X"D0", X"16", X"A6", X"D6", X"F0", X"37", X"C6", X"D6", X"A5", X"D3", X"38", X"E9", 
		X"28", X"90", X"04", X"85", X"D3", X"10", X"2A", X"20", X"6C", X"E5", X"D0", X"25", X"C9", X"12", X"D0", X"04", 
		X"A9", X"00", X"85", X"C7", X"C9", X"1D", X"D0", X"12", X"98", X"F0", X"09", X"20", X"A1", X"E8", X"88", X"84", 
		X"D3", X"4C", X"A8", X"E6", X"20", X"01", X"E7", X"4C", X"A8", X"E6", X"C9", X"13", X"D0", X"06", X"20", X"44", 
		X"E5", X"4C", X"A8", X"E6", X"09", X"80", X"20", X"CB", X"E8", X"4C", X"4F", X"EC", X"46", X"C9", X"A6", X"D6", 
		X"E8", X"E0", X"19", X"D0", X"03", X"20", X"EA", X"E8", X"B5", X"D9", X"10", X"F4", X"86", X"D6", X"4C", X"6C", 
		X"E5", X"A2", X"00", X"86", X"D8", X"86", X"C7", X"86", X"D4", X"86", X"D3", X"20", X"7C", X"E8", X"4C", X"A8", 
		X"E6", X"A2", X"02", X"A9", X"00", X"C5", X"D3", X"F0", X"07", X"18", X"69", X"28", X"CA", X"D0", X"F6", X"60", 
		X"C6", X"D6", X"60", X"A2", X"02", X"A9", X"27", X"C5", X"D3", X"F0", X"07", X"18", X"69", X"28", X"CA", X"D0", 
		X"F6", X"60", X"A6", X"D6", X"E0", X"19", X"F0", X"02", X"E6", X"D6", X"60", X"A2", X"0F", X"DD", X"DA", X"E8", 
		X"F0", X"04", X"CA", X"10", X"F8", X"60", X"8E", X"86", X"02", X"60", X"90", X"05", X"1C", X"9F", X"9C", X"1E", 
		X"1F", X"9E", X"81", X"95", X"96", X"97", X"98", X"99", X"9A", X"9B", X"A5", X"AC", X"48", X"A5", X"AD", X"48", 
		X"A5", X"AE", X"48", X"A5", X"AF", X"48", X"A2", X"FF", X"C6", X"D6", X"C6", X"C9", X"CE", X"A5", X"02", X"E8", 
		X"20", X"F0", X"E9", X"E0", X"18", X"B0", X"0C", X"BD", X"F1", X"EC", X"85", X"AC", X"B5", X"DA", X"20", X"C8", 
		X"E9", X"30", X"EC", X"20", X"FF", X"E9", X"A2", X"00", X"B5", X"D9", X"29", X"7F", X"B4", X"DA", X"10", X"02", 
		X"09", X"80", X"95", X"D9", X"E8", X"E0", X"18", X"D0", X"EF", X"A5", X"F1", X"09", X"80", X"85", X"F1", X"A5", 
		X"D9", X"10", X"C3", X"E6", X"D6", X"EE", X"A5", X"02", X"A9", X"7F", X"8D", X"00", X"DC", X"AD", X"01", X"DC", 
		X"C9", X"FB", X"08", X"A9", X"7F", X"8D", X"00", X"DC", X"28", X"D0", X"0B", X"A0", X"00", X"EA", X"CA", X"D0", 
		X"FC", X"88", X"D0", X"F9", X"84", X"C6", X"A6", X"D6", X"68", X"85", X"AF", X"68", X"85", X"AE", X"68", X"85", 
		X"AD", X"68", X"85", X"AC", X"60", X"A6", X"D6", X"E8", X"B5", X"D9", X"10", X"FB", X"8E", X"A5", X"02", X"E0", 
		X"18", X"F0", X"0E", X"90", X"0C", X"20", X"EA", X"E8", X"AE", X"A5", X"02", X"CA", X"C6", X"D6", X"4C", X"DA", 
		X"E6", X"A5", X"AC", X"48", X"A5", X"AD", X"48", X"A5", X"AE", X"48", X"A5", X"AF", X"48", X"A2", X"19", X"CA", 
		X"20", X"F0", X"E9", X"EC", X"A5", X"02", X"90", X"0E", X"F0", X"0C", X"BD", X"EF", X"EC", X"85", X"AC", X"B5", 
		X"D8", X"20", X"C8", X"E9", X"30", X"E9", X"20", X"FF", X"E9", X"A2", X"17", X"EC", X"A5", X"02", X"90", X"0F", 
		X"B5", X"DA", X"29", X"7F", X"B4", X"D9", X"10", X"02", X"09", X"80", X"95", X"DA", X"CA", X"D0", X"EC", X"AE", 
		X"A5", X"02", X"20", X"DA", X"E6", X"4C", X"58", X"E9", X"29", X"03", X"0D", X"88", X"02", X"85", X"AD", X"20", 
		X"E0", X"E9", X"A0", X"27", X"B1", X"AC", X"91", X"D1", X"B1", X"AE", X"91", X"F3", X"88", X"10", X"F5", X"60", 
		X"20", X"24", X"EA", X"A5", X"AC", X"85", X"AE", X"A5", X"AD", X"29", X"03", X"09", X"D8", X"85", X"AF", X"60", 
		X"BD", X"F0", X"EC", X"85", X"D1", X"B5", X"D9", X"29", X"03", X"0D", X"88", X"02", X"85", X"D2", X"60", X"A0", 
		X"27", X"20", X"F0", X"E9", X"20", X"24", X"EA", X"20", X"DA", X"E4", X"A9", X"20", X"91", X"D1", X"88", X"10", 
		X"F6", X"60", X"EA", X"A8", X"A9", X"02", X"85", X"CD", X"20", X"24", X"EA", X"98", X"A4", X"D3", X"91", X"D1", 
		X"8A", X"91", X"F3", X"60", X"A5", X"D1", X"85", X"F3", X"A5", X"D2", X"29", X"03", X"09", X"D8", X"85", X"F4", 
		X"60", X"20", X"EA", X"FF", X"A5", X"CC", X"D0", X"29", X"C6", X"CD", X"D0", X"25", X"A9", X"14", X"85", X"CD", 
		X"A4", X"D3", X"46", X"CF", X"AE", X"87", X"02", X"B1", X"D1", X"B0", X"11", X"E6", X"CF", X"85", X"CE", X"20", 
		X"24", X"EA", X"B1", X"F3", X"8D", X"87", X"02", X"AE", X"86", X"02", X"A5", X"CE", X"49", X"80", X"20", X"1C", 
		X"EA", X"A5", X"01", X"29", X"10", X"F0", X"0A", X"A0", X"00", X"84", X"C0", X"A5", X"01", X"09", X"20", X"D0", 
		X"08", X"A5", X"C0", X"D0", X"06", X"A5", X"01", X"29", X"1F", X"85", X"01", X"20", X"87", X"EA", X"AD", X"0D", 
		X"DC", X"68", X"A8", X"68", X"AA", X"68", X"40", X"A9", X"00", X"8D", X"8D", X"02", X"A0", X"40", X"84", X"CB", 
		X"8D", X"00", X"DC", X"AE", X"01", X"DC", X"E0", X"FF", X"F0", X"61", X"A8", X"A9", X"81", X"85", X"F5", X"A9", 
		X"EB", X"85", X"F6", X"A9", X"FE", X"8D", X"00", X"DC", X"A2", X"08", X"48", X"AD", X"01", X"DC", X"CD", X"01", 
		X"DC", X"D0", X"F8", X"4A", X"B0", X"16", X"48", X"B1", X"F5", X"C9", X"05", X"B0", X"0C", X"C9", X"03", X"F0", 
		X"08", X"0D", X"8D", X"02", X"8D", X"8D", X"02", X"10", X"02", X"84", X"CB", X"68", X"C8", X"C0", X"41", X"B0", 
		X"0B", X"CA", X"D0", X"DF", X"38", X"68", X"2A", X"8D", X"00", X"DC", X"D0", X"CC", X"68", X"6C", X"8F", X"02", 
		X"A4", X"CB", X"B1", X"F5", X"AA", X"C4", X"C5", X"F0", X"07", X"A0", X"10", X"8C", X"8C", X"02", X"D0", X"36", 
		X"29", X"7F", X"2C", X"8A", X"02", X"30", X"16", X"70", X"49", X"C9", X"7F", X"F0", X"29", X"C9", X"14", X"F0", 
		X"0C", X"C9", X"20", X"F0", X"08", X"C9", X"1D", X"F0", X"04", X"C9", X"11", X"D0", X"35", X"AC", X"8C", X"02", 
		X"F0", X"05", X"CE", X"8C", X"02", X"D0", X"2B", X"CE", X"8B", X"02", X"D0", X"26", X"A0", X"04", X"8C", X"8B", 
		X"02", X"A4", X"C6", X"88", X"10", X"1C", X"A4", X"CB", X"84", X"C5", X"AC", X"8D", X"02", X"8C", X"8E", X"02", 
		X"E0", X"FF", X"F0", X"0E", X"8A", X"A6", X"C6", X"EC", X"89", X"02", X"B0", X"06", X"9D", X"77", X"02", X"E8", 
		X"86", X"C6", X"A9", X"7F", X"8D", X"00", X"DC", X"60", X"AD", X"8D", X"02", X"C9", X"03", X"D0", X"15", X"CD", 
		X"8E", X"02", X"F0", X"EE", X"AD", X"91", X"02", X"30", X"1D", X"AD", X"18", X"D0", X"49", X"02", X"8D", X"18", 
		X"D0", X"4C", X"76", X"EB", X"0A", X"C9", X"08", X"90", X"02", X"A9", X"06", X"AA", X"BD", X"79", X"EB", X"85", 
		X"F5", X"BD", X"7A", X"EB", X"85", X"F6", X"4C", X"E0", X"EA", X"81", X"EB", X"C2", X"EB", X"03", X"EC", X"78", 
		X"EC", X"14", X"0D", X"1D", X"88", X"85", X"86", X"87", X"11", X"33", X"57", X"41", X"34", X"5A", X"53", X"45", 
		X"01", X"35", X"52", X"44", X"36", X"43", X"46", X"54", X"58", X"37", X"59", X"47", X"38", X"42", X"48", X"55", 
		X"56", X"39", X"49", X"4A", X"30", X"4D", X"4B", X"4F", X"4E", X"2B", X"50", X"4C", X"2D", X"2E", X"3A", X"40", 
		X"2C", X"5C", X"2A", X"3B", X"13", X"01", X"3D", X"5E", X"2F", X"31", X"5F", X"04", X"32", X"20", X"02", X"51", 
		X"03", X"FF", X"94", X"8D", X"9D", X"8C", X"89", X"8A", X"8B", X"91", X"23", X"D7", X"C1", X"24", X"DA", X"D3", 
		X"C5", X"01", X"25", X"D2", X"C4", X"26", X"C3", X"C6", X"D4", X"D8", X"27", X"D9", X"C7", X"28", X"C2", X"C8", 
		X"D5", X"D6", X"29", X"C9", X"CA", X"30", X"CD", X"CB", X"CF", X"CE", X"DB", X"D0", X"CC", X"DD", X"3E", X"5B", 
		X"BA", X"3C", X"A9", X"C0", X"5D", X"93", X"01", X"3D", X"DE", X"3F", X"21", X"5F", X"04", X"22", X"A0", X"02", 
		X"D1", X"83", X"FF", X"94", X"8D", X"9D", X"8C", X"89", X"8A", X"8B", X"91", X"96", X"B3", X"B0", X"97", X"AD", 
		X"AE", X"B1", X"01", X"98", X"B2", X"AC", X"99", X"BC", X"BB", X"A3", X"BD", X"9A", X"B7", X"A5", X"9B", X"BF", 
		X"B4", X"B8", X"BE", X"29", X"A2", X"B5", X"30", X"A7", X"A1", X"B9", X"AA", X"A6", X"AF", X"B6", X"DC", X"3E", 
		X"5B", X"A4", X"3C", X"A8", X"DF", X"5D", X"93", X"01", X"3D", X"DE", X"3F", X"81", X"5F", X"04", X"95", X"A0", 
		X"02", X"AB", X"83", X"FF", X"C9", X"0E", X"D0", X"07", X"AD", X"18", X"D0", X"09", X"02", X"D0", X"09", X"C9", 
		X"8E", X"D0", X"0B", X"AD", X"18", X"D0", X"29", X"FD", X"8D", X"18", X"D0", X"4C", X"A8", X"E6", X"C9", X"08", 
		X"D0", X"07", X"A9", X"80", X"0D", X"91", X"02", X"30", X"09", X"C9", X"09", X"D0", X"EE", X"A9", X"7F", X"2D", 
		X"91", X"02", X"8D", X"91", X"02", X"4C", X"A8", X"E6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
		X"1C", X"17", X"01", X"9F", X"1A", X"13", X"05", X"FF", X"9C", X"12", X"04", X"1E", X"03", X"06", X"14", X"18", 
		X"1F", X"19", X"07", X"9E", X"02", X"08", X"15", X"16", X"12", X"09", X"0A", X"92", X"0D", X"0B", X"0F", X"0E", 
		X"FF", X"10", X"0C", X"FF", X"FF", X"1B", X"00", X"FF", X"1C", X"FF", X"1D", X"FF", X"FF", X"1F", X"1E", X"FF", 
		X"90", X"06", X"FF", X"05", X"FF", X"FF", X"11", X"FF", X"FF", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"37", X"00", X"00", X"00", X"08", 
		X"00", X"14", X"0F", X"00", X"00", X"00", X"00", X"00", X"00", X"0E", X"06", X"01", X"02", X"03", X"04", X"00", 
		X"01", X"02", X"03", X"04", X"05", X"06", X"07", X"4C", X"4F", X"41", X"44", X"0D", X"52", X"55", X"4E", X"0D", 
		X"00", X"28", X"50", X"78", X"A0", X"C8", X"F0", X"18", X"40", X"68", X"90", X"B8", X"E0", X"08", X"30", X"58", 
		X"80", X"A8", X"D0", X"F8", X"20", X"48", X"70", X"98", X"C0", X"09", X"40", X"2C", X"09", X"20", X"20", X"A4", 
		X"F0", X"48", X"24", X"94", X"10", X"0A", X"38", X"66", X"A3", X"20", X"40", X"ED", X"46", X"94", X"46", X"A3", 
		X"68", X"85", X"95", X"78", X"20", X"97", X"EE", X"C9", X"3F", X"D0", X"03", X"20", X"85", X"EE", X"AD", X"00", 
		X"DD", X"09", X"08", X"8D", X"00", X"DD", X"78", X"20", X"8E", X"EE", X"20", X"97", X"EE", X"20", X"B3", X"EE", 
		X"78", X"20", X"97", X"EE", X"20", X"A9", X"EE", X"B0", X"64", X"20", X"85", X"EE", X"24", X"A3", X"10", X"0A", 
		X"20", X"A9", X"EE", X"90", X"FB", X"20", X"A9", X"EE", X"B0", X"FB", X"20", X"A9", X"EE", X"90", X"FB", X"20", 
		X"8E", X"EE", X"A9", X"08", X"85", X"A5", X"AD", X"00", X"DD", X"CD", X"00", X"DD", X"D0", X"F8", X"0A", X"90", 
		X"3F", X"66", X"95", X"B0", X"05", X"20", X"A0", X"EE", X"D0", X"03", X"20", X"97", X"EE", X"20", X"85", X"EE", 
		X"EA", X"EA", X"EA", X"EA", X"AD", X"00", X"DD", X"29", X"DF", X"09", X"10", X"8D", X"00", X"DD", X"C6", X"A5", 
		X"D0", X"D4", X"A9", X"04", X"8D", X"07", X"DC", X"A9", X"19", X"8D", X"0F", X"DC", X"AD", X"0D", X"DC", X"AD", 
		X"0D", X"DC", X"29", X"02", X"D0", X"0A", X"20", X"A9", X"EE", X"B0", X"F4", X"58", X"60", X"A9", X"80", X"2C", 
		X"A9", X"03", X"20", X"1C", X"FE", X"58", X"18", X"90", X"4A", X"85", X"95", X"20", X"36", X"ED", X"AD", X"00", 
		X"DD", X"29", X"F7", X"8D", X"00", X"DD", X"60", X"85", X"95", X"20", X"36", X"ED", X"78", X"20", X"A0", X"EE", 
		X"20", X"BE", X"ED", X"20", X"85", X"EE", X"20", X"A9", X"EE", X"30", X"FB", X"58", X"60", X"24", X"94", X"30", 
		X"05", X"38", X"66", X"94", X"D0", X"05", X"48", X"20", X"40", X"ED", X"68", X"85", X"95", X"18", X"60", X"78", 
		X"20", X"8E", X"EE", X"AD", X"00", X"DD", X"09", X"08", X"8D", X"00", X"DD", X"A9", X"5F", X"2C", X"A9", X"3F", 
		X"20", X"11", X"ED", X"20", X"BE", X"ED", X"8A", X"A2", X"0A", X"CA", X"D0", X"FD", X"AA", X"20", X"85", X"EE", 
		X"4C", X"97", X"EE", X"78", X"A9", X"00", X"85", X"A5", X"20", X"85", X"EE", X"20", X"A9", X"EE", X"10", X"FB", 
		X"A9", X"01", X"8D", X"07", X"DC", X"A9", X"19", X"8D", X"0F", X"DC", X"20", X"97", X"EE", X"AD", X"0D", X"DC", 
		X"AD", X"0D", X"DC", X"29", X"02", X"D0", X"07", X"20", X"A9", X"EE", X"30", X"F4", X"10", X"18", X"A5", X"A5", 
		X"F0", X"05", X"A9", X"02", X"4C", X"B2", X"ED", X"20", X"A0", X"EE", X"20", X"85", X"EE", X"A9", X"40", X"20", 
		X"1C", X"FE", X"E6", X"A5", X"D0", X"CA", X"A9", X"08", X"85", X"A5", X"AD", X"00", X"DD", X"CD", X"00", X"DD", 
		X"D0", X"F8", X"0A", X"10", X"F5", X"66", X"A4", X"AD", X"00", X"DD", X"CD", X"00", X"DD", X"D0", X"F8", X"0A", 
		X"30", X"F5", X"C6", X"A5", X"D0", X"E4", X"20", X"A0", X"EE", X"24", X"90", X"50", X"03", X"20", X"06", X"EE", 
		X"A5", X"A4", X"58", X"18", X"60", X"AD", X"00", X"DD", X"29", X"EF", X"8D", X"00", X"DD", X"60", X"AD", X"00", 
		X"DD", X"09", X"10", X"8D", X"00", X"DD", X"60", X"AD", X"00", X"DD", X"29", X"DF", X"8D", X"00", X"DD", X"60", 
		X"AD", X"00", X"DD", X"09", X"20", X"8D", X"00", X"DD", X"60", X"AD", X"00", X"DD", X"CD", X"00", X"DD", X"D0", 
		X"F8", X"0A", X"60", X"8A", X"A2", X"B8", X"CA", X"D0", X"FD", X"AA", X"60", X"A5", X"B4", X"F0", X"47", X"30", 
		X"3F", X"46", X"B6", X"A2", X"00", X"90", X"01", X"CA", X"8A", X"45", X"BD", X"85", X"BD", X"C6", X"B4", X"F0", 
		X"06", X"8A", X"29", X"04", X"85", X"B5", X"60", X"A9", X"20", X"2C", X"94", X"02", X"F0", X"14", X"30", X"1C", 
		X"70", X"14", X"A5", X"BD", X"D0", X"01", X"CA", X"C6", X"B4", X"AD", X"93", X"02", X"10", X"E3", X"C6", X"B4", 
		X"D0", X"DF", X"E6", X"B4", X"D0", X"F0", X"A5", X"BD", X"F0", X"ED", X"D0", X"EA", X"70", X"E9", X"50", X"E6", 
		X"E6", X"B4", X"A2", X"FF", X"D0", X"CB", X"AD", X"94", X"02", X"4A", X"90", X"07", X"2C", X"01", X"DD", X"10", 
		X"1D", X"50", X"1E", X"A9", X"00", X"85", X"BD", X"85", X"B5", X"AE", X"98", X"02", X"86", X"B4", X"AC", X"9D", 
		X"02", X"CC", X"9E", X"02", X"F0", X"13", X"B1", X"F9", X"85", X"B6", X"EE", X"9D", X"02", X"60", X"A9", X"40", 
		X"2C", X"A9", X"10", X"0D", X"97", X"02", X"8D", X"97", X"02", X"A9", X"01", X"8D", X"0D", X"DD", X"4D", X"A1", 
		X"02", X"09", X"80", X"8D", X"A1", X"02", X"8D", X"0D", X"DD", X"60", X"A2", X"09", X"A9", X"20", X"2C", X"93", 
		X"02", X"F0", X"01", X"CA", X"50", X"02", X"CA", X"CA", X"60", X"A6", X"A9", X"D0", X"33", X"C6", X"A8", X"F0", 
		X"36", X"30", X"0D", X"A5", X"A7", X"45", X"AB", X"85", X"AB", X"46", X"A7", X"66", X"AA", X"60", X"C6", X"A8", 
		X"A5", X"A7", X"F0", X"67", X"AD", X"93", X"02", X"0A", X"A9", X"01", X"65", X"A8", X"D0", X"EF", X"A9", X"90", 
		X"8D", X"0D", X"DD", X"0D", X"A1", X"02", X"8D", X"A1", X"02", X"85", X"A9", X"A9", X"02", X"4C", X"3B", X"EF", 
		X"A5", X"A7", X"D0", X"EA", X"4C", X"D3", X"E4", X"AC", X"9B", X"02", X"C8", X"CC", X"9C", X"02", X"F0", X"2A", 
		X"8C", X"9B", X"02", X"88", X"A5", X"AA", X"AE", X"98", X"02", X"E0", X"09", X"F0", X"04", X"4A", X"E8", X"D0", 
		X"F8", X"91", X"F7", X"A9", X"20", X"2C", X"94", X"02", X"F0", X"B4", X"30", X"B1", X"A5", X"A7", X"45", X"AB", 
		X"F0", X"03", X"70", X"A9", X"2C", X"50", X"A6", X"A9", X"01", X"2C", X"A9", X"04", X"2C", X"A9", X"80", X"2C", 
		X"A9", X"02", X"0D", X"97", X"02", X"8D", X"97", X"02", X"4C", X"7E", X"EF", X"A5", X"AA", X"D0", X"F1", X"F0", 
		X"EC", X"85", X"9A", X"AD", X"94", X"02", X"4A", X"90", X"29", X"A9", X"02", X"2C", X"01", X"DD", X"10", X"1D", 
		X"D0", X"20", X"AD", X"A1", X"02", X"29", X"02", X"D0", X"F9", X"2C", X"01", X"DD", X"70", X"FB", X"AD", X"01", 
		X"DD", X"09", X"02", X"8D", X"01", X"DD", X"2C", X"01", X"DD", X"70", X"07", X"30", X"F9", X"A9", X"40", X"8D", 
		X"97", X"02", X"18", X"60", X"20", X"28", X"F0", X"AC", X"9E", X"02", X"C8", X"CC", X"9D", X"02", X"F0", X"F4", 
		X"8C", X"9E", X"02", X"88", X"A5", X"9E", X"91", X"F9", X"AD", X"A1", X"02", X"4A", X"B0", X"1E", X"A9", X"10", 
		X"8D", X"0E", X"DD", X"AD", X"99", X"02", X"8D", X"04", X"DD", X"AD", X"9A", X"02", X"8D", X"05", X"DD", X"A9", 
		X"81", X"20", X"3B", X"EF", X"20", X"06", X"EF", X"A9", X"11", X"8D", X"0E", X"DD", X"60", X"85", X"99", X"AD", 
		X"94", X"02", X"4A", X"90", X"28", X"29", X"08", X"F0", X"24", X"A9", X"02", X"2C", X"01", X"DD", X"10", X"AD", 
		X"F0", X"22", X"AD", X"A1", X"02", X"4A", X"B0", X"FA", X"AD", X"01", X"DD", X"29", X"FD", X"8D", X"01", X"DD", 
		X"AD", X"01", X"DD", X"29", X"04", X"F0", X"F9", X"A9", X"90", X"18", X"4C", X"3B", X"EF", X"AD", X"A1", X"02", 
		X"29", X"12", X"F0", X"F3", X"18", X"60", X"AD", X"97", X"02", X"AC", X"9C", X"02", X"CC", X"9B", X"02", X"F0", 
		X"0B", X"29", X"F7", X"8D", X"97", X"02", X"B1", X"F7", X"EE", X"9C", X"02", X"60", X"09", X"08", X"8D", X"97", 
		X"02", X"A9", X"00", X"60", X"48", X"AD", X"A1", X"02", X"F0", X"11", X"AD", X"A1", X"02", X"29", X"03", X"D0", 
		X"F9", X"A9", X"10", X"8D", X"0D", X"DD", X"A9", X"00", X"8D", X"A1", X"02", X"68", X"60", X"0D", X"49", X"2F", 
		X"4F", X"20", X"45", X"52", X"52", X"4F", X"52", X"20", X"A3", X"0D", X"53", X"45", X"41", X"52", X"43", X"48", 
		X"49", X"4E", X"47", X"A0", X"46", X"4F", X"52", X"A0", X"0D", X"50", X"52", X"45", X"53", X"53", X"20", X"50", 
		X"4C", X"41", X"59", X"20", X"4F", X"4E", X"20", X"54", X"41", X"50", X"C5", X"50", X"52", X"45", X"53", X"53", 
		X"20", X"52", X"45", X"43", X"4F", X"52", X"44", X"20", X"26", X"20", X"50", X"4C", X"41", X"59", X"20", X"4F", 
		X"4E", X"20", X"54", X"41", X"50", X"C5", X"0D", X"4C", X"4F", X"41", X"44", X"49", X"4E", X"C7", X"0D", X"53", 
		X"41", X"56", X"49", X"4E", X"47", X"A0", X"0D", X"56", X"45", X"52", X"49", X"46", X"59", X"49", X"4E", X"C7", 
		X"0D", X"46", X"4F", X"55", X"4E", X"44", X"A0", X"0D", X"4F", X"4B", X"8D", X"24", X"9D", X"10", X"0D", X"B9", 
		X"BD", X"F0", X"08", X"29", X"7F", X"20", X"D2", X"FF", X"C8", X"28", X"10", X"F3", X"18", X"60", X"A5", X"99", 
		X"D0", X"08", X"A5", X"C6", X"F0", X"0F", X"78", X"4C", X"B4", X"E5", X"C9", X"02", X"D0", X"18", X"84", X"97", 
		X"20", X"86", X"F0", X"A4", X"97", X"18", X"60", X"A5", X"99", X"D0", X"0B", X"A5", X"D3", X"85", X"CA", X"A5", 
		X"D6", X"85", X"C9", X"4C", X"32", X"E6", X"C9", X"03", X"D0", X"09", X"85", X"D0", X"A5", X"D5", X"85", X"C8", 
		X"4C", X"32", X"E6", X"B0", X"38", X"C9", X"02", X"F0", X"3F", X"86", X"97", X"20", X"99", X"F1", X"B0", X"16", 
		X"48", X"20", X"99", X"F1", X"B0", X"0D", X"D0", X"05", X"A9", X"40", X"20", X"1C", X"FE", X"C6", X"A6", X"A6", 
		X"97", X"68", X"60", X"AA", X"68", X"8A", X"A6", X"97", X"60", X"20", X"0D", X"F8", X"D0", X"0B", X"20", X"41", 
		X"F8", X"B0", X"11", X"A9", X"00", X"85", X"A6", X"F0", X"F0", X"B1", X"B2", X"18", X"60", X"A5", X"90", X"F0", 
		X"04", X"A9", X"0D", X"18", X"60", X"4C", X"13", X"EE", X"20", X"4E", X"F1", X"B0", X"F7", X"C9", X"00", X"D0", 
		X"F2", X"AD", X"97", X"02", X"29", X"60", X"D0", X"E9", X"F0", X"EE", X"48", X"A5", X"9A", X"C9", X"03", X"D0", 
		X"04", X"68", X"4C", X"16", X"E7", X"90", X"04", X"68", X"4C", X"DD", X"ED", X"4A", X"68", X"85", X"9E", X"8A", 
		X"48", X"98", X"48", X"90", X"23", X"20", X"0D", X"F8", X"D0", X"0E", X"20", X"64", X"F8", X"B0", X"0E", X"A9", 
		X"02", X"A0", X"00", X"91", X"B2", X"C8", X"84", X"A6", X"A5", X"9E", X"91", X"B2", X"18", X"68", X"A8", X"68", 
		X"AA", X"A5", X"9E", X"90", X"02", X"A9", X"00", X"60", X"20", X"17", X"F0", X"4C", X"FC", X"F1", X"20", X"0F", 
		X"F3", X"F0", X"03", X"4C", X"01", X"F7", X"20", X"1F", X"F3", X"A5", X"BA", X"F0", X"16", X"C9", X"03", X"F0", 
		X"12", X"B0", X"14", X"C9", X"02", X"D0", X"03", X"4C", X"4D", X"F0", X"A6", X"B9", X"E0", X"60", X"F0", X"03", 
		X"4C", X"0A", X"F7", X"85", X"99", X"18", X"60", X"AA", X"20", X"09", X"ED", X"A5", X"B9", X"10", X"06", X"20", 
		X"CC", X"ED", X"4C", X"48", X"F2", X"20", X"C7", X"ED", X"8A", X"24", X"90", X"10", X"E6", X"4C", X"07", X"F7", 
		X"20", X"0F", X"F3", X"F0", X"03", X"4C", X"01", X"F7", X"20", X"1F", X"F3", X"A5", X"BA", X"D0", X"03", X"4C", 
		X"0D", X"F7", X"C9", X"03", X"F0", X"0F", X"B0", X"11", X"C9", X"02", X"D0", X"03", X"4C", X"E1", X"EF", X"A6", 
		X"B9", X"E0", X"60", X"F0", X"EA", X"85", X"9A", X"18", X"60", X"AA", X"20", X"0C", X"ED", X"A5", X"B9", X"10", 
		X"05", X"20", X"BE", X"ED", X"D0", X"03", X"20", X"B9", X"ED", X"8A", X"24", X"90", X"10", X"E7", X"4C", X"07", 
		X"F7", X"20", X"14", X"F3", X"F0", X"02", X"18", X"60", X"20", X"1F", X"F3", X"8A", X"48", X"A5", X"BA", X"F0", 
		X"50", X"C9", X"03", X"F0", X"4C", X"B0", X"47", X"C9", X"02", X"D0", X"1D", X"68", X"20", X"F2", X"F2", X"20", 
		X"83", X"F4", X"20", X"27", X"FE", X"A5", X"F8", X"F0", X"01", X"C8", X"A5", X"FA", X"F0", X"01", X"C8", X"A9", 
		X"00", X"85", X"F8", X"85", X"FA", X"4C", X"7D", X"F4", X"A5", X"B9", X"29", X"0F", X"F0", X"23", X"20", X"D0", 
		X"F7", X"A9", X"00", X"38", X"20", X"DD", X"F1", X"20", X"64", X"F8", X"90", X"04", X"68", X"A9", X"00", X"60", 
		X"A5", X"B9", X"C9", X"62", X"D0", X"0B", X"A9", X"05", X"20", X"6A", X"F7", X"4C", X"F1", X"F2", X"20", X"42", 
		X"F6", X"68", X"AA", X"C6", X"98", X"E4", X"98", X"F0", X"14", X"A4", X"98", X"B9", X"59", X"02", X"9D", X"59", 
		X"02", X"B9", X"63", X"02", X"9D", X"63", X"02", X"B9", X"6D", X"02", X"9D", X"6D", X"02", X"18", X"60", X"A9", 
		X"00", X"85", X"90", X"8A", X"A6", X"98", X"CA", X"30", X"15", X"DD", X"59", X"02", X"D0", X"F8", X"60", X"BD", 
		X"59", X"02", X"85", X"B8", X"BD", X"63", X"02", X"85", X"BA", X"BD", X"6D", X"02", X"85", X"B9", X"60", X"A9", 
		X"00", X"85", X"98", X"A2", X"03", X"E4", X"9A", X"B0", X"03", X"20", X"FE", X"ED", X"E4", X"99", X"B0", X"03", 
		X"20", X"EF", X"ED", X"86", X"9A", X"A9", X"00", X"85", X"99", X"60", X"A6", X"B8", X"D0", X"03", X"4C", X"0A", 
		X"F7", X"20", X"0F", X"F3", X"D0", X"03", X"4C", X"FE", X"F6", X"A6", X"98", X"E0", X"0A", X"90", X"03", X"4C", 
		X"FB", X"F6", X"E6", X"98", X"A5", X"B8", X"9D", X"59", X"02", X"A5", X"B9", X"09", X"60", X"85", X"B9", X"9D", 
		X"6D", X"02", X"A5", X"BA", X"9D", X"63", X"02", X"F0", X"5A", X"C9", X"03", X"F0", X"56", X"90", X"05", X"20", 
		X"D5", X"F3", X"90", X"4F", X"C9", X"02", X"D0", X"03", X"4C", X"09", X"F4", X"20", X"D0", X"F7", X"B0", X"03", 
		X"4C", X"13", X"F7", X"A5", X"B9", X"29", X"0F", X"D0", X"1F", X"20", X"17", X"F8", X"B0", X"36", X"20", X"AF", 
		X"F5", X"A5", X"B7", X"F0", X"0A", X"20", X"EA", X"F7", X"90", X"18", X"F0", X"28", X"4C", X"04", X"F7", X"20", 
		X"2C", X"F7", X"F0", X"20", X"90", X"0C", X"B0", X"F4", X"20", X"38", X"F8", X"B0", X"17", X"A9", X"04", X"20", 
		X"6A", X"F7", X"A9", X"BF", X"A4", X"B9", X"C0", X"60", X"F0", X"07", X"A0", X"00", X"A9", X"02", X"91", X"B2", 
		X"98", X"85", X"A6", X"18", X"60", X"A5", X"B9", X"30", X"FA", X"A4", X"B7", X"F0", X"F6", X"A9", X"00", X"85", 
		X"90", X"A5", X"BA", X"20", X"0C", X"ED", X"A5", X"B9", X"09", X"F0", X"20", X"B9", X"ED", X"A5", X"90", X"10", 
		X"05", X"68", X"68", X"4C", X"07", X"F7", X"A5", X"B7", X"F0", X"0C", X"A0", X"00", X"B1", X"BB", X"20", X"DD", 
		X"ED", X"C8", X"C4", X"B7", X"D0", X"F6", X"4C", X"54", X"F6", X"20", X"83", X"F4", X"8C", X"97", X"02", X"C4", 
		X"B7", X"F0", X"0A", X"B1", X"BB", X"99", X"93", X"02", X"C8", X"C0", X"04", X"D0", X"F2", X"20", X"4A", X"EF", 
		X"8E", X"98", X"02", X"AD", X"93", X"02", X"29", X"0F", X"F0", X"1C", X"0A", X"AA", X"AD", X"A6", X"02", X"D0", 
		X"09", X"BC", X"C1", X"FE", X"BD", X"C0", X"FE", X"4C", X"40", X"F4", X"BC", X"EB", X"E4", X"BD", X"EA", X"E4", 
		X"8C", X"96", X"02", X"8D", X"95", X"02", X"AD", X"95", X"02", X"0A", X"20", X"2E", X"FF", X"AD", X"94", X"02", 
		X"4A", X"90", X"09", X"AD", X"01", X"DD", X"0A", X"B0", X"03", X"20", X"0D", X"F0", X"AD", X"9B", X"02", X"8D", 
		X"9C", X"02", X"AD", X"9E", X"02", X"8D", X"9D", X"02", X"20", X"27", X"FE", X"A5", X"F8", X"D0", X"05", X"88", 
		X"84", X"F8", X"86", X"F7", X"A5", X"FA", X"D0", X"05", X"88", X"84", X"FA", X"86", X"F9", X"38", X"A9", X"F0", 
		X"4C", X"2D", X"FE", X"A9", X"7F", X"8D", X"0D", X"DD", X"A9", X"06", X"8D", X"03", X"DD", X"8D", X"01", X"DD", 
		X"A9", X"04", X"0D", X"00", X"DD", X"8D", X"00", X"DD", X"A0", X"00", X"8C", X"A1", X"02", X"60", X"86", X"C3", 
		X"84", X"C4", X"6C", X"30", X"03", X"85", X"93", X"A9", X"00", X"85", X"90", X"A5", X"BA", X"D0", X"03", X"4C", 
		X"13", X"F7", X"C9", X"03", X"F0", X"F9", X"90", X"7B", X"A4", X"B7", X"D0", X"03", X"4C", X"10", X"F7", X"A6", 
		X"B9", X"20", X"AF", X"F5", X"A9", X"60", X"85", X"B9", X"20", X"D5", X"F3", X"A5", X"BA", X"20", X"09", X"ED", 
		X"A5", X"B9", X"20", X"C7", X"ED", X"20", X"13", X"EE", X"85", X"AE", X"A5", X"90", X"4A", X"4A", X"B0", X"50", 
		X"20", X"13", X"EE", X"85", X"AF", X"8A", X"D0", X"08", X"A5", X"C3", X"85", X"AE", X"A5", X"C4", X"85", X"AF", 
		X"20", X"D2", X"F5", X"A9", X"FD", X"25", X"90", X"85", X"90", X"20", X"E1", X"FF", X"D0", X"03", X"4C", X"33", 
		X"F6", X"20", X"13", X"EE", X"AA", X"A5", X"90", X"4A", X"4A", X"B0", X"E8", X"8A", X"A4", X"93", X"F0", X"0C", 
		X"A0", X"00", X"D1", X"AE", X"F0", X"08", X"A9", X"10", X"20", X"1C", X"FE", X"2C", X"91", X"AE", X"E6", X"AE", 
		X"D0", X"02", X"E6", X"AF", X"24", X"90", X"50", X"CB", X"20", X"EF", X"ED", X"20", X"42", X"F6", X"90", X"79", 
		X"4C", X"04", X"F7", X"4A", X"B0", X"03", X"4C", X"13", X"F7", X"20", X"D0", X"F7", X"B0", X"03", X"4C", X"13", 
		X"F7", X"20", X"17", X"F8", X"B0", X"68", X"20", X"AF", X"F5", X"A5", X"B7", X"F0", X"09", X"20", X"EA", X"F7", 
		X"90", X"0B", X"F0", X"5A", X"B0", X"DA", X"20", X"2C", X"F7", X"F0", X"53", X"B0", X"D3", X"A5", X"90", X"29", 
		X"10", X"38", X"D0", X"4A", X"E0", X"01", X"F0", X"11", X"E0", X"03", X"D0", X"DD", X"A0", X"01", X"B1", X"B2", 
		X"85", X"C3", X"C8", X"B1", X"B2", X"85", X"C4", X"B0", X"04", X"A5", X"B9", X"D0", X"EF", X"A0", X"03", X"B1", 
		X"B2", X"A0", X"01", X"F1", X"B2", X"AA", X"A0", X"04", X"B1", X"B2", X"A0", X"02", X"F1", X"B2", X"A8", X"18", 
		X"8A", X"65", X"C3", X"85", X"AE", X"98", X"65", X"C4", X"85", X"AF", X"A5", X"C3", X"85", X"C1", X"A5", X"C4", 
		X"85", X"C2", X"20", X"D2", X"F5", X"20", X"4A", X"F8", X"24", X"18", X"A6", X"AE", X"A4", X"AF", X"60", X"A5", 
		X"9D", X"10", X"1E", X"A0", X"0C", X"20", X"2F", X"F1", X"A5", X"B7", X"F0", X"15", X"A0", X"17", X"20", X"2F", 
		X"F1", X"A4", X"B7", X"F0", X"0C", X"A0", X"00", X"B1", X"BB", X"20", X"D2", X"FF", X"C8", X"C4", X"B7", X"D0", 
		X"F6", X"60", X"A0", X"49", X"A5", X"93", X"F0", X"02", X"A0", X"59", X"4C", X"2B", X"F1", X"86", X"AE", X"84", 
		X"AF", X"AA", X"B5", X"00", X"85", X"C1", X"B5", X"01", X"85", X"C2", X"6C", X"32", X"03", X"A5", X"BA", X"D0", 
		X"03", X"4C", X"13", X"F7", X"C9", X"03", X"F0", X"F9", X"90", X"5F", X"A9", X"61", X"85", X"B9", X"A4", X"B7", 
		X"D0", X"03", X"4C", X"10", X"F7", X"20", X"D5", X"F3", X"20", X"8F", X"F6", X"A5", X"BA", X"20", X"0C", X"ED", 
		X"A5", X"B9", X"20", X"B9", X"ED", X"A0", X"00", X"20", X"8E", X"FB", X"A5", X"AC", X"20", X"DD", X"ED", X"A5", 
		X"AD", X"20", X"DD", X"ED", X"20", X"D1", X"FC", X"B0", X"16", X"B1", X"AC", X"20", X"DD", X"ED", X"20", X"E1", 
		X"FF", X"D0", X"07", X"20", X"42", X"F6", X"A9", X"00", X"38", X"60", X"20", X"DB", X"FC", X"D0", X"E5", X"20", 
		X"FE", X"ED", X"24", X"B9", X"30", X"11", X"A5", X"BA", X"20", X"0C", X"ED", X"A5", X"B9", X"29", X"EF", X"09", 
		X"E0", X"20", X"B9", X"ED", X"20", X"FE", X"ED", X"18", X"60", X"4A", X"B0", X"03", X"4C", X"13", X"F7", X"20", 
		X"D0", X"F7", X"90", X"8D", X"20", X"38", X"F8", X"B0", X"25", X"20", X"8F", X"F6", X"A2", X"03", X"A5", X"B9", 
		X"29", X"01", X"D0", X"02", X"A2", X"01", X"8A", X"20", X"6A", X"F7", X"B0", X"12", X"20", X"67", X"F8", X"B0", 
		X"0D", X"A5", X"B9", X"29", X"02", X"F0", X"06", X"A9", X"05", X"20", X"6A", X"F7", X"24", X"18", X"60", X"A5", 
		X"9D", X"10", X"FB", X"A0", X"51", X"20", X"2F", X"F1", X"4C", X"C1", X"F5", X"A2", X"00", X"E6", X"A2", X"D0", 
		X"06", X"E6", X"A1", X"D0", X"02", X"E6", X"A0", X"38", X"A5", X"A2", X"E9", X"01", X"A5", X"A1", X"E9", X"1A", 
		X"A5", X"A0", X"E9", X"4F", X"90", X"06", X"86", X"A0", X"86", X"A1", X"86", X"A2", X"AD", X"01", X"DC", X"CD", 
		X"01", X"DC", X"D0", X"F8", X"AA", X"30", X"13", X"A2", X"BD", X"8E", X"00", X"DC", X"AE", X"01", X"DC", X"EC", 
		X"01", X"DC", X"D0", X"F8", X"8D", X"00", X"DC", X"E8", X"D0", X"02", X"85", X"91", X"60", X"78", X"A5", X"A2", 
		X"A6", X"A1", X"A4", X"A0", X"78", X"85", X"A2", X"86", X"A1", X"84", X"A0", X"58", X"60", X"A5", X"91", X"C9", 
		X"7F", X"D0", X"07", X"08", X"20", X"CC", X"FF", X"85", X"C6", X"28", X"60", X"A9", X"01", X"2C", X"A9", X"02", 
		X"2C", X"A9", X"03", X"2C", X"A9", X"04", X"2C", X"A9", X"05", X"2C", X"A9", X"06", X"2C", X"A9", X"07", X"2C", 
		X"A9", X"08", X"2C", X"A9", X"09", X"48", X"20", X"CC", X"FF", X"A0", X"00", X"24", X"9D", X"50", X"0A", X"20", 
		X"2F", X"F1", X"68", X"48", X"09", X"30", X"20", X"D2", X"FF", X"68", X"38", X"60", X"A5", X"93", X"48", X"20", 
		X"41", X"F8", X"68", X"85", X"93", X"B0", X"32", X"A0", X"00", X"B1", X"B2", X"C9", X"05", X"F0", X"2A", X"C9", 
		X"01", X"F0", X"08", X"C9", X"03", X"F0", X"04", X"C9", X"04", X"D0", X"E1", X"AA", X"24", X"9D", X"10", X"17", 
		X"A0", X"63", X"20", X"2F", X"F1", X"A0", X"05", X"B1", X"B2", X"20", X"D2", X"FF", X"C8", X"C0", X"15", X"D0", 
		X"F6", X"A5", X"A1", X"20", X"E0", X"E4", X"EA", X"18", X"88", X"60", X"85", X"9E", X"20", X"D0", X"F7", X"90", 
		X"5E", X"A5", X"C2", X"48", X"A5", X"C1", X"48", X"A5", X"AF", X"48", X"A5", X"AE", X"48", X"A0", X"BF", X"A9", 
		X"20", X"91", X"B2", X"88", X"D0", X"FB", X"A5", X"9E", X"91", X"B2", X"C8", X"A5", X"C1", X"91", X"B2", X"C8", 
		X"A5", X"C2", X"91", X"B2", X"C8", X"A5", X"AE", X"91", X"B2", X"C8", X"A5", X"AF", X"91", X"B2", X"C8", X"84", 
		X"9F", X"A0", X"00", X"84", X"9E", X"A4", X"9E", X"C4", X"B7", X"F0", X"0C", X"B1", X"BB", X"A4", X"9F", X"91", 
		X"B2", X"E6", X"9E", X"E6", X"9F", X"D0", X"EE", X"20", X"D7", X"F7", X"A9", X"69", X"85", X"AB", X"20", X"6B", 
		X"F8", X"A8", X"68", X"85", X"AE", X"68", X"85", X"AF", X"68", X"85", X"C1", X"68", X"85", X"C2", X"98", X"60", 
		X"A6", X"B2", X"A4", X"B3", X"C0", X"02", X"60", X"20", X"D0", X"F7", X"8A", X"85", X"C1", X"18", X"69", X"C0", 
		X"85", X"AE", X"98", X"85", X"C2", X"69", X"00", X"85", X"AF", X"60", X"20", X"2C", X"F7", X"B0", X"1D", X"A0", 
		X"05", X"84", X"9F", X"A0", X"00", X"84", X"9E", X"C4", X"B7", X"F0", X"10", X"B1", X"BB", X"A4", X"9F", X"D1", 
		X"B2", X"D0", X"E7", X"E6", X"9E", X"E6", X"9F", X"A4", X"9E", X"D0", X"EC", X"18", X"60", X"20", X"D0", X"F7", 
		X"E6", X"A6", X"A4", X"A6", X"C0", X"C0", X"60", X"20", X"2E", X"F8", X"F0", X"1A", X"A0", X"1B", X"20", X"2F", 
		X"F1", X"20", X"D0", X"F8", X"20", X"2E", X"F8", X"D0", X"F8", X"A0", X"6A", X"4C", X"2F", X"F1", X"A9", X"10", 
		X"24", X"01", X"D0", X"02", X"24", X"01", X"18", X"60", X"20", X"2E", X"F8", X"F0", X"F9", X"A0", X"2E", X"D0", 
		X"DD", X"A9", X"00", X"85", X"90", X"85", X"93", X"20", X"D7", X"F7", X"20", X"17", X"F8", X"B0", X"1F", X"78", 
		X"A9", X"00", X"85", X"AA", X"85", X"B4", X"85", X"B0", X"85", X"9E", X"85", X"9F", X"85", X"9C", X"A9", X"90", 
		X"A2", X"0E", X"D0", X"11", X"20", X"D7", X"F7", X"A9", X"14", X"85", X"AB", X"20", X"38", X"F8", X"B0", X"6C", 
		X"78", X"A9", X"82", X"A2", X"08", X"A0", X"7F", X"8C", X"0D", X"DC", X"8D", X"0D", X"DC", X"AD", X"0E", X"DC", 
		X"09", X"19", X"8D", X"0F", X"DC", X"29", X"91", X"8D", X"A2", X"02", X"20", X"A4", X"F0", X"AD", X"11", X"D0", 
		X"29", X"EF", X"8D", X"11", X"D0", X"AD", X"14", X"03", X"8D", X"9F", X"02", X"AD", X"15", X"03", X"8D", X"A0", 
		X"02", X"20", X"BD", X"FC", X"A9", X"02", X"85", X"BE", X"20", X"97", X"FB", X"A5", X"01", X"29", X"1F", X"85", 
		X"01", X"85", X"C0", X"A2", X"FF", X"A0", X"FF", X"88", X"D0", X"FD", X"CA", X"D0", X"F8", X"58", X"AD", X"A0", 
		X"02", X"CD", X"15", X"03", X"18", X"F0", X"15", X"20", X"D0", X"F8", X"20", X"BC", X"F6", X"4C", X"BE", X"F8", 
		X"20", X"E1", X"FF", X"18", X"D0", X"0B", X"20", X"93", X"FC", X"38", X"68", X"68", X"A9", X"00", X"8D", X"A0", 
		X"02", X"60", X"86", X"B1", X"A5", X"B0", X"0A", X"0A", X"18", X"65", X"B0", X"18", X"65", X"B1", X"85", X"B1", 
		X"A9", X"00", X"24", X"B0", X"30", X"01", X"2A", X"06", X"B1", X"2A", X"06", X"B1", X"2A", X"AA", X"AD", X"06", 
		X"DC", X"C9", X"16", X"90", X"F9", X"65", X"B1", X"8D", X"04", X"DC", X"8A", X"6D", X"07", X"DC", X"8D", X"05", 
		X"DC", X"AD", X"A2", X"02", X"8D", X"0E", X"DC", X"8D", X"A4", X"02", X"AD", X"0D", X"DC", X"29", X"10", X"F0", 
		X"09", X"A9", X"F9", X"48", X"A9", X"2A", X"48", X"4C", X"43", X"FF", X"58", X"60", X"AE", X"07", X"DC", X"A0", 
		X"FF", X"98", X"ED", X"06", X"DC", X"EC", X"07", X"DC", X"D0", X"F2", X"86", X"B1", X"AA", X"8C", X"06", X"DC", 
		X"8C", X"07", X"DC", X"A9", X"19", X"8D", X"0F", X"DC", X"AD", X"0D", X"DC", X"8D", X"A3", X"02", X"98", X"E5", 
		X"B1", X"86", X"B1", X"4A", X"66", X"B1", X"4A", X"66", X"B1", X"A5", X"B0", X"18", X"69", X"3C", X"C5", X"B1", 
		X"B0", X"4A", X"A6", X"9C", X"F0", X"03", X"4C", X"60", X"FA", X"A6", X"A3", X"30", X"1B", X"A2", X"00", X"69", 
		X"30", X"65", X"B0", X"C5", X"B1", X"B0", X"1C", X"E8", X"69", X"26", X"65", X"B0", X"C5", X"B1", X"B0", X"17", 
		X"69", X"2C", X"65", X"B0", X"C5", X"B1", X"90", X"03", X"4C", X"10", X"FA", X"A5", X"B4", X"F0", X"1D", X"85", 
		X"A8", X"D0", X"19", X"E6", X"A9", X"B0", X"02", X"C6", X"A9", X"38", X"E9", X"13", X"E5", X"B1", X"65", X"92", 
		X"85", X"92", X"A5", X"A4", X"49", X"01", X"85", X"A4", X"F0", X"2B", X"86", X"D7", X"A5", X"B4", X"F0", X"22", 
		X"AD", X"A3", X"02", X"29", X"01", X"D0", X"05", X"AD", X"A4", X"02", X"D0", X"16", X"A9", X"00", X"85", X"A4", 
		X"8D", X"A4", X"02", X"A5", X"A3", X"10", X"30", X"30", X"BF", X"A2", X"A6", X"20", X"E2", X"F8", X"A5", X"9B", 
		X"D0", X"B9", X"4C", X"BC", X"FE", X"A5", X"92", X"F0", X"07", X"30", X"03", X"C6", X"B0", X"2C", X"E6", X"B0", 
		X"A9", X"00", X"85", X"92", X"E4", X"D7", X"D0", X"0F", X"8A", X"D0", X"A0", X"A5", X"A9", X"30", X"BD", X"C9", 
		X"10", X"90", X"B9", X"85", X"96", X"B0", X"B5", X"8A", X"45", X"9B", X"85", X"9B", X"A5", X"B4", X"F0", X"D2", 
		X"C6", X"A3", X"30", X"C5", X"46", X"D7", X"66", X"BF", X"A2", X"DA", X"20", X"E2", X"F8", X"4C", X"BC", X"FE", 
		X"A5", X"96", X"F0", X"04", X"A5", X"B4", X"F0", X"07", X"A5", X"A3", X"30", X"03", X"4C", X"97", X"F9", X"46", 
		X"B1", X"A9", X"93", X"38", X"E5", X"B1", X"65", X"B0", X"0A", X"AA", X"20", X"E2", X"F8", X"E6", X"9C", X"A5", 
		X"B4", X"D0", X"11", X"A5", X"96", X"F0", X"26", X"85", X"A8", X"A9", X"00", X"85", X"96", X"A9", X"81", X"8D", 
		X"0D", X"DC", X"85", X"B4", X"A5", X"96", X"85", X"B5", X"F0", X"09", X"A9", X"00", X"85", X"B4", X"A9", X"01", 
		X"8D", X"0D", X"DC", X"A5", X"BF", X"85", X"BD", X"A5", X"A8", X"05", X"A9", X"85", X"B6", X"4C", X"BC", X"FE", 
		X"20", X"97", X"FB", X"85", X"9C", X"A2", X"DA", X"20", X"E2", X"F8", X"A5", X"BE", X"F0", X"02", X"85", X"A7", 
		X"A9", X"0F", X"24", X"AA", X"10", X"17", X"A5", X"B5", X"D0", X"0C", X"A6", X"BE", X"CA", X"D0", X"0B", X"A9", 
		X"08", X"20", X"1C", X"FE", X"D0", X"04", X"A9", X"00", X"85", X"AA", X"4C", X"BC", X"FE", X"70", X"31", X"D0", 
		X"18", X"A5", X"B5", X"D0", X"F5", X"A5", X"B6", X"D0", X"F1", X"A5", X"A7", X"4A", X"A5", X"BD", X"30", X"03", 
		X"90", X"18", X"18", X"B0", X"15", X"29", X"0F", X"85", X"AA", X"C6", X"AA", X"D0", X"DD", X"A9", X"40", X"85", 
		X"AA", X"20", X"8E", X"FB", X"A9", X"00", X"85", X"AB", X"F0", X"D0", X"A9", X"80", X"85", X"AA", X"D0", X"CA", 
		X"A5", X"B5", X"F0", X"0A", X"A9", X"04", X"20", X"1C", X"FE", X"A9", X"00", X"4C", X"4A", X"FB", X"20", X"D1", 
		X"FC", X"90", X"03", X"4C", X"48", X"FB", X"A6", X"A7", X"CA", X"F0", X"2D", X"A5", X"93", X"F0", X"0C", X"A0", 
		X"00", X"A5", X"BD", X"D1", X"AC", X"F0", X"04", X"A9", X"01", X"85", X"B6", X"A5", X"B6", X"F0", X"4B", X"A2", 
		X"3D", X"E4", X"9E", X"90", X"3E", X"A6", X"9E", X"A5", X"AD", X"9D", X"01", X"01", X"A5", X"AC", X"9D", X"00", 
		X"01", X"E8", X"E8", X"86", X"9E", X"4C", X"3A", X"FB", X"A6", X"9F", X"E4", X"9E", X"F0", X"35", X"A5", X"AC", 
		X"DD", X"00", X"01", X"D0", X"2E", X"A5", X"AD", X"DD", X"01", X"01", X"D0", X"27", X"E6", X"9F", X"E6", X"9F", 
		X"A5", X"93", X"F0", X"0B", X"A5", X"BD", X"A0", X"00", X"D1", X"AC", X"F0", X"17", X"C8", X"84", X"B6", X"A5", 
		X"B6", X"F0", X"07", X"A9", X"10", X"20", X"1C", X"FE", X"D0", X"09", X"A5", X"93", X"D0", X"05", X"A8", X"A5", 
		X"BD", X"91", X"AC", X"20", X"DB", X"FC", X"D0", X"43", X"A9", X"80", X"85", X"AA", X"78", X"A2", X"01", X"8E", 
		X"0D", X"DC", X"AE", X"0D", X"DC", X"A6", X"BE", X"CA", X"30", X"02", X"86", X"BE", X"C6", X"A7", X"F0", X"08", 
		X"A5", X"9E", X"D0", X"27", X"85", X"BE", X"F0", X"23", X"20", X"93", X"FC", X"20", X"8E", X"FB", X"A0", X"00", 
		X"84", X"AB", X"B1", X"AC", X"45", X"AB", X"85", X"AB", X"20", X"DB", X"FC", X"20", X"D1", X"FC", X"90", X"F2", 
		X"A5", X"AB", X"45", X"BD", X"F0", X"05", X"A9", X"20", X"20", X"1C", X"FE", X"4C", X"BC", X"FE", X"A5", X"C2", 
		X"85", X"AD", X"A5", X"C1", X"85", X"AC", X"60", X"A9", X"08", X"85", X"A3", X"A9", X"00", X"85", X"A4", X"85", 
		X"A8", X"85", X"9B", X"85", X"A9", X"60", X"A5", X"BD", X"4A", X"A9", X"60", X"90", X"02", X"A9", X"B0", X"A2", 
		X"00", X"8D", X"06", X"DC", X"8E", X"07", X"DC", X"AD", X"0D", X"DC", X"A9", X"19", X"8D", X"0F", X"DC", X"A5", 
		X"01", X"49", X"08", X"85", X"01", X"29", X"08", X"60", X"38", X"66", X"B6", X"30", X"3C", X"A5", X"A8", X"D0", 
		X"12", X"A9", X"10", X"A2", X"01", X"20", X"B1", X"FB", X"D0", X"2F", X"E6", X"A8", X"A5", X"B6", X"10", X"29", 
		X"4C", X"57", X"FC", X"A5", X"A9", X"D0", X"09", X"20", X"AD", X"FB", X"D0", X"1D", X"E6", X"A9", X"D0", X"19", 
		X"20", X"A6", X"FB", X"D0", X"14", X"A5", X"A4", X"49", X"01", X"85", X"A4", X"F0", X"0F", X"A5", X"BD", X"49", 
		X"01", X"85", X"BD", X"29", X"01", X"45", X"9B", X"85", X"9B", X"4C", X"BC", X"FE", X"46", X"BD", X"C6", X"A3", 
		X"A5", X"A3", X"F0", X"3A", X"10", X"F3", X"20", X"97", X"FB", X"58", X"A5", X"A5", X"F0", X"12", X"A2", X"00", 
		X"86", X"D7", X"C6", X"A5", X"A6", X"BE", X"E0", X"02", X"D0", X"02", X"09", X"80", X"85", X"BD", X"D0", X"D9", 
		X"20", X"D1", X"FC", X"90", X"0A", X"D0", X"91", X"E6", X"AD", X"A5", X"D7", X"85", X"BD", X"B0", X"CA", X"A0", 
		X"00", X"B1", X"AC", X"85", X"BD", X"45", X"D7", X"85", X"D7", X"20", X"DB", X"FC", X"D0", X"BB", X"A5", X"9B", 
		X"49", X"01", X"85", X"BD", X"4C", X"BC", X"FE", X"C6", X"BE", X"D0", X"03", X"20", X"CA", X"FC", X"A9", X"50", 
		X"85", X"A7", X"A2", X"08", X"78", X"20", X"BD", X"FC", X"D0", X"EA", X"A9", X"78", X"20", X"AF", X"FB", X"D0", 
		X"E3", X"C6", X"A7", X"D0", X"DF", X"20", X"97", X"FB", X"C6", X"AB", X"10", X"D8", X"A2", X"0A", X"20", X"BD", 
		X"FC", X"58", X"E6", X"AB", X"A5", X"BE", X"F0", X"30", X"20", X"8E", X"FB", X"A2", X"09", X"86", X"A5", X"86", 
		X"B6", X"D0", X"83", X"08", X"78", X"AD", X"11", X"D0", X"09", X"10", X"8D", X"11", X"D0", X"20", X"CA", X"FC", 
		X"A9", X"7F", X"8D", X"0D", X"DC", X"20", X"DD", X"FD", X"AD", X"A0", X"02", X"F0", X"09", X"8D", X"15", X"03", 
		X"AD", X"9F", X"02", X"8D", X"14", X"03", X"28", X"60", X"20", X"93", X"FC", X"F0", X"97", X"BD", X"93", X"FD", 
		X"8D", X"14", X"03", X"BD", X"94", X"FD", X"8D", X"15", X"03", X"60", X"A5", X"01", X"09", X"20", X"85", X"01", 
		X"60", X"38", X"A5", X"AC", X"E5", X"AE", X"A5", X"AD", X"E5", X"AF", X"60", X"E6", X"AC", X"D0", X"02", X"E6", 
		X"AD", X"60", X"A2", X"FF", X"78", X"9A", X"D8", X"20", X"02", X"FD", X"D0", X"03", X"6C", X"00", X"80", X"8E", 
		X"16", X"D0", X"20", X"A3", X"FD", X"20", X"50", X"FD", X"20", X"15", X"FD", X"20", X"5B", X"FF", X"58", X"6C", 
		X"00", X"A0", X"A2", X"05", X"BD", X"0F", X"FD", X"DD", X"03", X"80", X"D0", X"03", X"CA", X"D0", X"F5", X"60", 
		X"C3", X"C2", X"CD", X"38", X"30", X"A2", X"30", X"A0", X"FD", X"18", X"86", X"C3", X"84", X"C4", X"A0", X"1F", 
		X"B9", X"14", X"03", X"B0", X"02", X"B1", X"C3", X"91", X"C3", X"99", X"14", X"03", X"88", X"10", X"F1", X"60", 
		X"31", X"EA", X"66", X"FE", X"47", X"FE", X"4A", X"F3", X"91", X"F2", X"0E", X"F2", X"50", X"F2", X"33", X"F3", 
		X"57", X"F1", X"CA", X"F1", X"ED", X"F6", X"3E", X"F1", X"2F", X"F3", X"66", X"FE", X"A5", X"F4", X"ED", X"F5", 
		X"A9", X"00", X"A8", X"99", X"02", X"00", X"99", X"00", X"02", X"99", X"00", X"03", X"C8", X"D0", X"F4", X"A2", 
		X"3C", X"A0", X"03", X"86", X"B2", X"84", X"B3", X"A8", X"A9", X"03", X"85", X"C2", X"E6", X"C2", X"B1", X"C1", 
		X"AA", X"A9", X"55", X"91", X"C1", X"D1", X"C1", X"D0", X"0F", X"2A", X"91", X"C1", X"D1", X"C1", X"D0", X"08", 
		X"8A", X"91", X"C1", X"C8", X"D0", X"E8", X"F0", X"E4", X"98", X"AA", X"A4", X"C2", X"18", X"20", X"2D", X"FE", 
		X"A9", X"08", X"8D", X"82", X"02", X"A9", X"04", X"8D", X"88", X"02", X"60", X"6A", X"FC", X"CD", X"FB", X"31", 
		X"EA", X"2C", X"F9", X"A9", X"7F", X"8D", X"0D", X"DC", X"8D", X"0D", X"DD", X"8D", X"00", X"DC", X"A9", X"08", 
		X"8D", X"0E", X"DC", X"8D", X"0E", X"DD", X"8D", X"0F", X"DC", X"8D", X"0F", X"DD", X"A2", X"00", X"8E", X"03", 
		X"DC", X"8E", X"03", X"DD", X"8E", X"18", X"D4", X"CA", X"8E", X"02", X"DC", X"A9", X"07", X"8D", X"00", X"DD", 
		X"A9", X"3F", X"8D", X"02", X"DD", X"A9", X"E7", X"85", X"01", X"A9", X"2F", X"85", X"00", X"AD", X"A6", X"02", 
		X"F0", X"0A", X"A9", X"25", X"8D", X"04", X"DC", X"A9", X"40", X"4C", X"F3", X"FD", X"A9", X"95", X"8D", X"04", 
		X"DC", X"A9", X"42", X"8D", X"05", X"DC", X"4C", X"6E", X"FF", X"85", X"B7", X"86", X"BB", X"84", X"BC", X"60", 
		X"85", X"B8", X"86", X"BA", X"84", X"B9", X"60", X"A5", X"BA", X"C9", X"02", X"D0", X"0D", X"AD", X"97", X"02", 
		X"48", X"A9", X"00", X"8D", X"97", X"02", X"68", X"60", X"85", X"9D", X"A5", X"90", X"05", X"90", X"85", X"90", 
		X"60", X"8D", X"85", X"02", X"60", X"90", X"06", X"AE", X"83", X"02", X"AC", X"84", X"02", X"8E", X"83", X"02", 
		X"8C", X"84", X"02", X"60", X"90", X"06", X"AE", X"81", X"02", X"AC", X"82", X"02", X"8E", X"81", X"02", X"8C", 
		X"82", X"02", X"60", X"78", X"6C", X"18", X"03", X"48", X"8A", X"48", X"98", X"48", X"A9", X"7F", X"8D", X"0D", 
		X"DD", X"AC", X"0D", X"DD", X"30", X"1C", X"20", X"02", X"FD", X"D0", X"03", X"6C", X"02", X"80", X"20", X"BC", 
		X"F6", X"20", X"E1", X"FF", X"D0", X"0C", X"20", X"15", X"FD", X"20", X"A3", X"FD", X"20", X"18", X"E5", X"6C", 
		X"02", X"A0", X"98", X"2D", X"A1", X"02", X"AA", X"29", X"01", X"F0", X"28", X"AD", X"00", X"DD", X"29", X"FB", 
		X"05", X"B5", X"8D", X"00", X"DD", X"AD", X"A1", X"02", X"8D", X"0D", X"DD", X"8A", X"29", X"12", X"F0", X"0D", 
		X"29", X"02", X"F0", X"06", X"20", X"D6", X"FE", X"4C", X"9D", X"FE", X"20", X"07", X"FF", X"20", X"BB", X"EE", 
		X"4C", X"B6", X"FE", X"8A", X"29", X"02", X"F0", X"06", X"20", X"D6", X"FE", X"4C", X"B6", X"FE", X"8A", X"29", 
		X"10", X"F0", X"03", X"20", X"07", X"FF", X"AD", X"A1", X"02", X"8D", X"0D", X"DD", X"68", X"A8", X"68", X"AA", 
		X"68", X"40", X"C1", X"27", X"3E", X"1A", X"C5", X"11", X"74", X"0E", X"ED", X"0C", X"45", X"06", X"F0", X"02", 
		X"46", X"01", X"B8", X"00", X"71", X"00", X"AD", X"01", X"DD", X"29", X"01", X"85", X"A7", X"AD", X"06", X"DD", 
		X"E9", X"1C", X"6D", X"99", X"02", X"8D", X"06", X"DD", X"AD", X"07", X"DD", X"6D", X"9A", X"02", X"8D", X"07", 
		X"DD", X"A9", X"11", X"8D", X"0F", X"DD", X"AD", X"A1", X"02", X"8D", X"0D", X"DD", X"A9", X"FF", X"8D", X"06", 
		X"DD", X"8D", X"07", X"DD", X"4C", X"59", X"EF", X"AD", X"95", X"02", X"8D", X"06", X"DD", X"AD", X"96", X"02", 
		X"8D", X"07", X"DD", X"A9", X"11", X"8D", X"0F", X"DD", X"A9", X"12", X"4D", X"A1", X"02", X"8D", X"A1", X"02", 
		X"A9", X"FF", X"8D", X"06", X"DD", X"8D", X"07", X"DD", X"AE", X"98", X"02", X"86", X"A8", X"60", X"AA", X"AD", 
		X"96", X"02", X"2A", X"A8", X"8A", X"69", X"C8", X"8D", X"99", X"02", X"98", X"69", X"00", X"8D", X"9A", X"02", 
		X"60", X"EA", X"EA", X"08", X"68", X"29", X"EF", X"48", X"48", X"8A", X"48", X"98", X"48", X"BA", X"BD", X"04", 
		X"01", X"29", X"10", X"F0", X"03", X"6C", X"16", X"03", X"6C", X"14", X"03", X"20", X"18", X"E5", X"AD", X"12", 
		X"D0", X"D0", X"FB", X"AD", X"19", X"D0", X"29", X"01", X"8D", X"A6", X"02", X"4C", X"DD", X"FD", X"A9", X"81", 
		X"8D", X"0D", X"DC", X"AD", X"0E", X"DC", X"29", X"80", X"09", X"11", X"8D", X"0E", X"DC", X"4C", X"8E", X"EE", 
		X"03", X"4C", X"5B", X"FF", X"4C", X"A3", X"FD", X"4C", X"50", X"FD", X"4C", X"15", X"FD", X"4C", X"1A", X"FD", 
		X"4C", X"18", X"FE", X"4C", X"B9", X"ED", X"4C", X"C7", X"ED", X"4C", X"25", X"FE", X"4C", X"34", X"FE", X"4C", 
		X"87", X"EA", X"4C", X"21", X"FE", X"4C", X"13", X"EE", X"4C", X"DD", X"ED", X"4C", X"EF", X"ED", X"4C", X"FE", 
		X"ED", X"4C", X"0C", X"ED", X"4C", X"09", X"ED", X"4C", X"07", X"FE", X"4C", X"00", X"FE", X"4C", X"F9", X"FD", 
		X"6C", X"1A", X"03", X"6C", X"1C", X"03", X"6C", X"1E", X"03", X"6C", X"20", X"03", X"6C", X"22", X"03", X"6C", 
		X"24", X"03", X"6C", X"26", X"03", X"4C", X"9E", X"F4", X"4C", X"DD", X"F5", X"4C", X"E4", X"F6", X"4C", X"DD", 
		X"F6", X"6C", X"28", X"03", X"6C", X"2A", X"03", X"6C", X"2C", X"03", X"4C", X"9B", X"F6", X"4C", X"05", X"E5", 
		X"4C", X"0A", X"E5", X"4C", X"00", X"E5", X"52", X"52", X"42", X"59", X"43", X"FE", X"E2", X"FC", X"48", X"FF" 
	);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			do <= romData(to_integer(addr)) after 2 ns;
		end if;
	end process;
end architecture;

